////////////////////////////////////////////////////////////////////////////////
// 
// Company: {{COMPANY}}
// Author: {{AUTHOR}}
//
// Create Date: {{DATE}}
// Module Name: {{MODULE_NAME}}
// Description:
//     {{DESCRIPTION}}
//
////////////////////////////////////////////////////////////////////////////////

mon module